library IEEE;
use IEEE.std_logic_1164.all;

entity This is
    port (
        a: in STD_LOGIC_VECTOR (3 downto 0);
        b: in STD_LOGIC_VECTOR (3 downto 0);
        c: out STD_LOGIC_VECTOR (3 downto 0)
    );
end This;

architecture This_arch of This is
begin
  -- <<enter your statements here>>
end This_arch;
